module tft_pic
(
input wire tft_clk_9m , //输入工作时钟,频率9MHz
input wire sys_rst_n , //输入复位信号,低电平有效
input wire [9:0] pix_x , //输入有效显示区域像素点X轴坐标
input wire [9:0] pix_y , //输入有效显示区域像素点Y轴坐标
input wire  ageb_sig1 ,
input wire  ageb_sig2 ,
output reg [15:0] pix_data //输出像素点色彩信息

);
////
//\* Parameter and Internal Signal \//
////
parameter H_VALID = 10'd480 , //行有效数据
V_VALID = 10'd272 ; //场有效数据
parameter CHAR_B_H= 10'd112 , //字符开始X轴坐标
CHAR_B_V= 10'd104 ; //字符开始Y轴坐标
parameter CHAR_W = 10'd256 , //字符宽度
CHAR_H = 10'd64 ; //字符高度
parameter BLACK = 16'h0000, //黑色
GOLDEN = 16'hFEC0; //金色
//wire define
wire [9:0] char_x ; //字符显示X轴坐标
wire [9:0] char_y ; //字符显示Y轴坐标
//reg define
reg [255:0] char [63:0] ; //字符数据
////
//\* Main Code \//
////
//字符显示坐标
assign char_x = (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
&& ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
? (pix_x - CHAR_B_H) : 10'h3FF;
assign char_y = (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
&& ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
? (pix_y - CHAR_B_V) : 10'h3FF;
//char:字符数据
always@(posedge tft_clk_9m)
if (ageb_sig1 == 1'b1)
begin
char[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[3] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[4] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[5] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[6] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[7] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[8] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[9] <= 256'h0000000000000000000000010000000004000000003E00000000003000000000;
char[10] <= 256'h06000000000000000000000F800000001E000000003E0000000000F800000000;
char[11] <= 256'h0F8000000000000000000007C00000000F800000003E00000000007C00000000;
char[12] <= 256'h0FE00FFFFFFFE00000000003E000000007C00000003E00000000003E00000000;
char[13] <= 256'h07F00FFFFFFFE00000000001F000000003E00000003E00007FFFFFFFFFFFFF80;
char[14] <= 256'h01FC0FFFFFFFE00001FFFFFFFFFFFF8003F00000003E00007FFFFFFFFFFFFF80;
char[15] <= 256'h007F0F000001E00001FFFFFFFFFFFF8001F80000003E00007FFFFFFFFFFFFF80;
char[16] <= 256'h003E0F000001E00001FFFFFFFFFFFF8000F80000003E00000000000000000000;
char[17] <= 256'h00080F000001E00001E00000003C000000787FFFFFFFFF800000000000000000;
char[18] <= 256'h00000FFFFFFFE00001E00780003C000000207FFFFFFFFF80003FFFFFFFFE0000;
char[19] <= 256'h00000FFFFFFFE00001E00780003C000000007FFFFFFFFF80003FFFFFFFFE0000;
char[20] <= 256'h30000FFFFFFFE00001E00780003C000000000000003E0000003FFFFFFFFE0000;
char[21] <= 256'h7C000F000001E00001EFFFFFFFFFFF0000000000003E0000003C0000001E0000;
char[22] <= 256'hFF000F000001E00001EFFFFFFFFFFF0000000000003E0000003C0000001E0000;
char[23] <= 256'h3FC00F000001E00001EFFFFFFFFFFF007FF00200003E0000003C0000001E0000;
char[24] <= 256'h0FE00FFFFFFFE00001E00780003C00007FF00780003E0000003C0000001E0000;
char[25] <= 256'h03F80FFFFFFFE00001E00780003C00007FF007C0003E0000003FFFFFFFFE0000;
char[26] <= 256'h01F00FFFFFFFE00001E00780003C000000F003E0003E0000003FFFFFFFFE0000;
char[27] <= 256'h00400F000001E00001E00780003C000000F001F0003E0000003FFFFFFFFE0000;
char[28] <= 256'h00000F000001E00001E007FFFFFC000000F000F8003E0000003C0000001E0000;
char[29] <= 256'h000000000000000001E007FFFFFC000000F0007C003E00000000000000000000;
char[30] <= 256'h000000000000000001E007FFFFFC000000F0003E003E00000FFFFFFFFFFFFC00;
char[31] <= 256'h00007FFFFFFFF80001E00780003C000000F0001F803E00000FFFFFFFFFFFFC00;
char[32] <= 256'h01807FFFFFFFF80001E000000000000000F0000F003E00000FFFFFFFFFFFFC00;
char[33] <= 256'h01F07FFFFFFFF80001E000000000000000F00004003E00000F00000000003C00;
char[34] <= 256'h03F0780F03C0780001E3FFFFFFFFC00000F00000003E00000F00000000003C00;
char[35] <= 256'h03E0780F03C0780003E3FFFFFFFFC00000F00000003E00000F00000000003C00;
char[36] <= 256'h03E0780F03C0780003C3FFFFFFFFC00000F00000003E00000F00FFFFFFC03C00;
char[37] <= 256'h03E0780F03C0780003C01F00001F800000F00000003E00000F00FFFFFFC03C00;
char[38] <= 256'h07C0780F03C0780003C00FC0003F000000F00000007E00000F00FFFFFFC03C00;
char[39] <= 256'h07C0780F03C0780003C003F000FC000000F00003FFFC00000F00F00003C03C00;
char[40] <= 256'h07C0780F03C0780007C001FC03F0000001F00001FFF800000F00F00003C03C00;
char[41] <= 256'h0F80780F03C078000780007F1FE0000003F80001FFF000000F00F00003C03C00;
char[42] <= 256'h0F80780F03C078000F80003FFF8000000FFC0000000000000F00FFFFFFC03C00;
char[43] <= 256'h0F80780F03C078000F800007FC0000001F9F8000000000000F00FFFFFFC03C00;
char[44] <= 256'h1F0FFFFFFFFFFF801F00007FFF8000007F0FF800000000000F00FFFFFFC03C00;
char[45] <= 256'h1F0FFFFFFFFFFF801F0007FFFFF800003C07FFFFFFFFFF800F00F00000007C00;
char[46] <= 256'h1F0FFFFFFFFFFF803E01FFFC0FFFC0003800FFFFFFFFFF800F00000003FFF800;
char[47] <= 256'h3E000000000000007C7FFFC000FFFF80100007FFFFFFFF000F00000001FFF800;
char[48] <= 256'h06000000000000001C3FF800000FFF0000000000000000000F00000001FFE000;
char[49] <= 256'h0000000000000000081E000000001E0000000000000000000000000000000000;
char[50] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[51] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[52] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[53] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[54] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[55] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[56] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[57] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[58] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[59] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[60] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;

end
else if (ageb_sig2 == 1'b0 )
begin
char[0]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[1]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[2]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[3]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[4]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[5]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[6]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[7]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[8]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[9]  <= 256'h0000000000000000000000010000000004000000003E00000000003000000000;
char[10]  <= 256'h00000000000000000000000F800000001E000000003E0000000000F800000000;
char[11]  <= 256'h060000000000000000000007C00000000F800000003E00000000007C00000000;
char[12]  <= 256'h0F001FFFFFFFF00000000003E000000007C00000003E00000000003E00000000;
char[13]  <= 256'h0FC01FFFFFFFF00000000001F000000003E00000003E00007FFFFFFFFFFFFF80;
char[14]  <= 256'h07F01FFFFFFFF00001FFFFFFFFFFFF8003F00000003E00007FFFFFFFFFFFFF80;
char[15]  <= 256'h01F81E000000F00001FFFFFFFFFFFF8001F80000003E00007FFFFFFFFFFFFF80;
char[16]  <= 256'h00FE1E000000F00001FFFFFFFFFFFF8000F80000003E00000000000000000000;
char[17]  <= 256'h003C1E000000F00001E00000003C000000787FFFFFFFFF800000000000000000;
char[18]  <= 256'h00101FFFFFFFF00001E00780003C000000207FFFFFFFFF80003FFFFFFFFE0000;
char[19]  <= 256'h00001FFFFFFFF00001E00780003C000000007FFFFFFFFF80003FFFFFFFFE0000;
char[20]  <= 256'h00001FFFFFFFF00001E00780003C000000000000003E0000003FFFFFFFFE0000;
char[21]  <= 256'h18001E000000F00001EFFFFFFFFFFF0000000000003E0000003C0000001E0000;
char[22]  <= 256'h3E001E000000F00001EFFFFFFFFFFF0000000000003E0000003C0000001E0000;
char[23]  <= 256'h7F801E000000F00001EFFFFFFFFFFF007FF00200003E0000003C0000001E0000;
char[24]  <= 256'h1FE01FFFFFFFF00001E00780003C00007FF00780003E0000003C0000001E0000;
char[25]  <= 256'h07F81FFFFFFFF00001E00780003C00007FF007C0003E0000003FFFFFFFFE0000;
char[26]  <= 256'h01FC1FFFFFFFF00001E00780003C000000F003E0003E0000003FFFFFFFFE0000;
char[27]  <= 256'h00F81E000000F00001E00780003C000000F001F0003E0000003FFFFFFFFE0000;
char[28]  <= 256'h0020001E01E0000001E007FFFFFC000000F000F8003E0000003C0000001E0000;
char[29]  <= 256'h0000001E01E0000001E007FFFFFC000000F0007C003E00000000000000000000;
char[30]  <= 256'h0000001E01E0000001E007FFFFFC000000F0003E003E00000FFFFFFFFFFFFC00;
char[31]  <= 256'h0000301E01E0080001E00780003C000000F0001F803E00000FFFFFFFFFFFFC00;
char[32]  <= 256'h0180F81E01E01F0001E000000000000000F0000F003E00000FFFFFFFFFFFFC00;
char[33]  <= 256'h01F07C1E01E03E0001E000000000000000F00004003E00000F00000000003C00;
char[34]  <= 256'h03F07C1E01E07C0001E3FFFFFFFFC00000F00000003E00000F00000000003C00;
char[35]  <= 256'h03E03E1E01E07C0003E3FFFFFFFFC00000F00000003E00000F00000000003C00;
char[36]  <= 256'h03E01E1E01E0F80003C3FFFFFFFFC00000F00000003E00000F00FFFFFFC03C00;
char[37]  <= 256'h03E01F1E01E1F00003C01F00001F800000F00000003E00000F00FFFFFFC03C00;
char[38]  <= 256'h07C00F1E01E3E00003C00FC0003F000000F00000007E00000F00FFFFFFC03C00;
char[39]  <= 256'h07C00F9E01E7C00003C003F000FC000000F00003FFFC00000F00F00003C03C00;
char[40]  <= 256'h07C0041E01E0800007C001FC03F0000001F00001FFF800000F00F00003C03C00;
char[41]  <= 256'h0F80001E01E000000780007F1FE0000003F80001FFF000000F00F00003C03C00;
char[42]  <= 256'h0F80001E01E000000F80003FFF8000000FFC0000000000000F00FFFFFFC03C00;
char[43]  <= 256'h0F80001E01E000000F800007FC0000001F9F8000000000000F00FFFFFFC03C00;
char[44]  <= 256'h1F03FFFFFFFFFF001F00007FFF8000007F0FF800000000000F00FFFFFFC03C00;
char[45]  <= 256'h1F03FFFFFFFFFF001F0007FFFFF800003C07FFFFFFFFFF800F00F00000007C00;
char[46]  <= 256'h1F03FFFFFFFFFF003E01FFFC0FFFC0003800FFFFFFFFFF800F00000003FFF800;
char[47]  <= 256'h3E000000000000007C7FFFC000FFFF80100007FFFFFFFF000F00000001FFF800;
char[48]  <= 256'h06000000000000001C3FF800000FFF0000000000000000000F00000001FFE000;
char[49]  <= 256'h0000000000000000081E000000001E0000000000000000000000000000000000;
char[50]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[51]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[52]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[53]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[54]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[55]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[56]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[57]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[58]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[59]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[60]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[61]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[62]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[63]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;


end
//pix_data:输出像素点色彩信息,根据当前像素点坐标指定当前像素点颜色数据
always@(posedge tft_clk_9m or negedge sys_rst_n)
if(sys_rst_n == 1'b0)
pix_data <= BLACK;
else if(((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
&& ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
begin
if(char[char_y][10'd255 - char_x] == 1'b1)
pix_data <= GOLDEN;
else
pix_data <= BLACK;
end
else
pix_data <= BLACK;
endmodule